module mma1(clk,reset,w,x,u);
input clk,reset;
input signed [15:0] w[0:2][0:2];
input  signed [15:0] x[0:2][0:63];
output signed [31:0] u[0:2][0:63];



//1
wxpe block1(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][0],x[1][0],x[2][0],u[0][0],u[1][0],u[2][0]);

//2
wxpe block2(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][1],x[1][1],x[2][1],u[0][1],u[1][1],u[2][1]);

//3
wxpe block3(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][2],x[1][2],x[2][2],u[0][2],u[1][2],u[2][2]);

//4
wxpe block4(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][3],x[1][3],x[2][3],u[0][3],u[1][3],u[2][3]);


//5
wxpe block5(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][4],x[1][4],x[2][4],u[0][4],u[1][4],u[2][4]);


//6
wxpe block6(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][5],x[1][5],x[2][5],u[0][5],u[1][5],u[2][5]);

//7
wxpe block7(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][6],x[1][6],x[2][6],u[0][6],u[1][6],u[2][6]);


//8
wxpe block8(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][7],x[1][7],x[2][7],u[0][7],u[1][7],u[2][7]);



//9
wxpe block9(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][8],x[1][8],x[2][8],u[0][8],u[1][8],u[2][8]);


//10
wxpe block10(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][9],x[1][9],x[2][9],u[0][9],u[1][9],u[2][9]);


//11
wxpe block11(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][10],x[1][10],x[2][10],u[0][10],u[1][10],u[2][10]);


//12
wxpe block12(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][11],x[1][11],x[2][11],u[0][11],u[1][11],u[2][11]);


//13
wxpe block13(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][12],x[1][12],x[2][12],u[0][12],u[1][12],u[2][12]);


//14
wxpe block14(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][13],x[1][13],x[2][13],u[0][13],u[1][13],u[2][13]);


//15
wxpe block15(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][14],x[1][14],x[2][14],u[0][14],u[1][14],u[2][14]);


//16
wxpe block16(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][15],x[1][15],x[2][15],u[0][15],u[1][15],u[2][15]);


//17
wxpe block17(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][16],x[1][16],x[2][16],u[0][16],u[1][16],u[2][16]);



//18
wxpe block18(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][17],x[1][17],x[2][17],u[0][17],u[1][17],u[2][17]);


//19
wxpe block19(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][18],x[1][18],x[2][18],u[0][18],u[1][18],u[2][18]);


//20
wxpe block20(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][19],x[1][19],x[2][19],u[0][19],u[1][19],u[2][19]);


//21
wxpe block21(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][20],x[1][20],x[2][20],u[0][20],u[1][20],u[2][20]);

//22
wxpe block22(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][21],x[1][21],x[2][21],u[0][21],u[1][21],u[2][21]);


//23
wxpe block23(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][22],x[1][22],x[2][22],u[0][22],u[1][22],u[2][22]);





//24
wxpe block24(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][23],x[1][23],x[2][23],u[0][23],u[1][23],u[2][23]);

//25
wxpe block25(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][24],x[1][24],x[2][24],u[0][24],u[1][24],u[2][24]);


//26
wxpe block26(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][25],x[1][25],x[2][25],u[0][25],u[1][25],u[2][25]);



//27
wxpe block27(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][26],x[1][26],x[2][26],u[0][26],u[1][26],u[2][26]);


//28
wxpe block28(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][27],x[1][27],x[2][27],u[0][27],u[1][27],u[2][27]);


//29
wxpe block29(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][28],x[1][28],x[2][28],u[0][28],u[1][28],u[2][28]);


//30
wxpe block30(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][29],x[1][29],x[2][29],u[0][29],u[1][29],u[2][29]);


//31
wxpe block31(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][30],x[1][30],x[2][30],u[0][30],u[1][30],u[2][30]);


//32
wxpe block32(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][31],x[1][31],x[2][31],u[0][31],u[1][31],u[2][31]);

//33
wxpe block33(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][32],x[1][32],x[2][32],u[0][32],u[1][32],u[2][32]);



//34
wxpe block34(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][33],x[1][33],x[2][33],u[0][33],u[1][33],u[2][33]);


//35
wxpe block35(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][34],x[1][34],x[2][34],u[0][34],u[1][34],u[2][34]);


//36
wxpe block36(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][35],x[1][35],x[2][35],u[0][35],u[1][35],u[2][35]);


//37
wxpe block37(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][36],x[1][36],x[2][36],u[0][36],u[1][36],u[2][36]);



//38
wxpe block38(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][37],x[1][37],x[2][37],u[0][37],u[1][37],u[2][37]);


//39
wxpe block39(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][38],x[1][38],x[2][38],u[0][38],u[1][38],u[2][38]);

//40
wxpe block40(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][39],x[1][39],x[2][39],u[0][39],u[1][39],u[2][39]);


//41
wxpe block41(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][40],x[1][40],x[2][40],u[0][40],u[1][40],u[2][40]);


//42
wxpe block42(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][41],x[1][41],x[2][41],u[0][41],u[1][41],u[2][41]);


//43
wxpe block43(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][42],x[1][42],x[2][42],u[0][42],u[1][42],u[2][42]);

//44
wxpe block44(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][43],x[1][43],x[2][43],u[0][43],u[1][43],u[2][43]);


//45
wxpe block45(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][44],x[1][44],x[2][44],u[0][44],u[1][44],u[2][44]);


//46
wxpe block46(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][45],x[1][45],x[2][45],u[0][45],u[1][45],u[2][45]);

//47
wxpe block47(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][46],x[1][46],x[2][46],u[0][46],u[1][46],u[2][46]);


//48
wxpe block48(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][47],x[1][47],x[2][47],u[0][47],u[1][47],u[2][47]);


//49
wxpe block49(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][48],x[1][48],x[2][48],u[0][48],u[1][48],u[2][48]);


//50
wxpe block50(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][49],x[1][49],x[2][49],u[0][49],u[1][49],u[2][49]);


//51
wxpe block51(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][50],x[1][50],x[2][50],u[0][50],u[1][50],u[2][50]);


//52
wxpe block52(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][51],x[1][51],x[2][51],u[0][51],u[1][51],u[2][51]);


//53
wxpe block53(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][52],x[1][52],x[2][52],u[0][52],u[1][52],u[2][52]);


//54
wxpe block54(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][53],x[1][53],x[2][53],u[0][53],u[1][53],u[2][53]);


//55
wxpe block55(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][54],x[1][54],x[2][54],u[0][54],u[1][54],u[2][54]);


//56
wxpe block56(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][55],x[1][55],x[2][55],u[0][55],u[1][55],u[2][55]);


//57
wxpe block57(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][56],x[1][56],x[2][56],u[0][56],u[1][56],u[2][56]);



//58
wxpe block58(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][57],x[1][57],x[2][57],u[0][57],u[1][57],u[2][57]);


//59
wxpe block59(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][58],x[1][58],x[2][58],u[0][58],u[1][58],u[2][58]);



//60
wxpe block60(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][59],x[1][59],x[2][59],u[0][59],u[1][59],u[2][59]);

//61
wxpe block61(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][60],x[1][60],x[2][60],u[0][60],u[1][60],u[2][60]);


//62
wxpe block62(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][61],x[1][61],x[2][61],u[0][61],u[1][61],u[2][61]);


//63
wxpe block63(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][62],x[1][62],x[2][62],u[0][62],u[1][62],u[2][62]);


//64

wxpe block64(clk,reset,w[0][0],w[0][1],w[0][2],w[1][0],w[1][1],w[1][2],w[2][0],w[2][1],w[2][2],x[0][63],x[1][63],x[2][63],u[0][63],u[1][63],u[2][63]);


endmodule


